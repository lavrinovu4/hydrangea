`ifndef __GLOBAL_DEF__
`define __GLOBAL_DEF__

`define US 1_000
`define MS (1_000 * `US)
`define S (1_000 * `MS)

`endif  //!__GLOBAL_DEF__
