`ifndef __GLOBAL_DEFINE__
`define __GLOBAL_DEFINE__

`timescale 1ns/10ps

`define SQ_INC 0
`define SQ_JMP 1
`define SQ_LOOP 2


`endif  //!__GLOBAL_DEFINE__
