
class cache_data;

  bit  [29:0] cache_addr  = 0 ;
  bit         cache_req  = 0 ;
  bit [31:0]   cache_data  ;
  bit          cache_ack   ;

endclass : cache_data
